RL Circuit Transient Response
r1 va vb 1000
l1 vb 0 1
*piecewise linear input voltage
vin va 0 pwl (0 0 10ms 0 11ms 5v 20ms 5v)
*transient analysis for 20ms, step size 0.02ms
.tran 0.02ms 20ms
.control
run
hardcopy rl_transient_01.ps v(va) v(vb)
set height=99999
print v(va) v(vb) > tmp.txt
.endc
.end